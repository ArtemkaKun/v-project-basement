module main

fn main() {
	println('Hellow, vorld!')
}