module main

fn test_main() {
	println('Hello Vorld')
}
